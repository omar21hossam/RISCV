class lsu_master_sequencer #(
    type REQ = lsu_sequence_item,
    type RSP = REQ
) extends uvm_sequencer #(lsu_sequence_item);

  //==================================================================================
  // Registeration
  //==================================================================================
  `uvm_component_utils(lsu_master_sequencer)

  //==================================================================================
  // Function: Constructor
  //==================================================================================
  function new(string name = "lsu_master_sequencer", uvm_component parent = null);
    super.new(name, parent);
  endfunction

endclass
