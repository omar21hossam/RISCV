package classes_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh";
  `include "lsu_sequence_item.svh";
  `include "lsu_master_sequence.svh";
  `include "lsu_master_sequencer.svh";
  `include "lsu_master_driver.svh";
  `include "lsu_master_monitor.svh";
  `include "lsu_master_agent.svh";
  `include "lsu_slave_sequence.svh";
  `include "lsu_slave_sequencer.svh";
  `include "lsu_slave_driver.svh";
  `include "lsu_slave_monitor.svh";
  `include "lsu_slave_agent.svh";
  `include "lsu_subscriber.svh";
  `include "lsu_scoreboard.svh";
  `include "lsu_env.svh";
  `include "lsu_test.svh";
endpackage

