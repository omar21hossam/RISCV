`timescale 1ns/1ps  
`include "ALU_interface.svh"
module riscv_alu_top_tb(
);
//==============================================================================
// Description: Parameters
//==============================================================================
parameter ClkPeriod = 10;
//==============================================================================
// Description: Clock
//==============================================================================
bit           clk_tb;
//==============================================================================
// Description: Include the packages
//==============================================================================
import uvm_pkg::*;
import package_uvm::*;
//==============================================================================
//Description: Clock generator
//==============================================================================
initial begin:clk_gen
forever begin
#(ClkPeriod/2) clk_tb = ~ clk_tb;
end 
end
//==============================================================================
//Description: Interface
//==============================================================================
ALU_interface  intf1(clk_tb);
//==============================================================================
//Description: DUT
//==============================================================================
    

//==============================================================================
//Description: Main block
//==============================================================================
initial begin
uvm_config_db#(virtual ALU_interface)::set(null,"uvm_test_top","top2test",intf1);
run_test();		
end

//==============================================================================
// initial begin
//     $dumpfile("riscv_top_tb.vcd");
//     $dumpvars(0,riscv_alu_top_tb);
//     $display("Starting simulation");
// end

    
endmodule