package classes_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh";
  `include "lsu_sequence_item.svh";
  `include "lsu_sequence.svh";
  `include "lsu_sequencer.svh";
  `include "lsu_subscriber.svh";
  `include "lsu_scoreboard.svh";
  `include "lsu_driver.svh";
  `include "lsu_active_driver.svh";
  `include "lsu_monitor.svh";
  `include "lsu_agent.svh";
  `include "lsu_env.svh";
  `include "lsu_test.svh";
endpackage

