class riscv_config_obj extends uvm_object;

  //==================================================================================
  // Registeration
  //==================================================================================
  `uvm_object_utils(riscv_config_obj);



  //==================================================================================
  // Agent State Enum
  //==================================================================================
  uvm_active_passive_enum active;

  //==================================================================================
  // Function: Constructor
  //==================================================================================
  function new(string name = "riscv_config_obj");
    super.new(name);
  endfunction

endclass
