class mul_seq_item extends uvm_sequence_item;
  `uvm_object_utils(mul_seq_item)

  // Declare the data members
  

  // Constructor
  function new(string name = "mul_seq_item");
    super.new(name);
  endfunction

  // Print function for debugging
endclass : mul_seq_item