`define LSU_PATH DUT.core_i.load_store_unit
