class alu_seq_item extends uvm_sequence_item;
  `uvm_object_utils(alu_seq_item)

  // Declare the data members
  

  // Constructor
  function new(string name = "alu_seq_item");
    super.new(name);
  endfunction

  // Print function for debugging
endclass : alu_seq_item