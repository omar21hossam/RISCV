//include all the interfaces used in the testbench
`include "ALU_DIV/tb_files/ALU_interface.svh"
