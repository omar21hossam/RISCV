package riscv_pkg;
  typedef enum logic [6:0] {
    OPCODE_LUI    = 7'b0110111,  //  (55)  : LUI Instruction
    OPCODE_AUIPC  = 7'b0010111,  //  (23)  : AUIPC Instruction
    OPCODE_JAL    = 7'b1101111,  //  (111) : JAL Instruction
    OPCODE_JALR   = 7'b1100111,  //  (103) : JALR Instruction
    OPCODE_BRANCH = 7'b1100011,  //  (99)  : Branch Instructions
    OPCODE_LOAD   = 7'b0000011,  //  (3)   : Load instructions
    OPCODE_STORE  = 7'b0100011,  //  (35)  : Store Instructions
    OPCODE_OP_IMM = 7'b0010011,  //  (19)  : I-type instructions
    OPCODE_OP     = 7'b0110011   //  (51)  : R-type Instructions
  } opcode_e;

  typedef enum logic [2:0] {
    ADD_SUB = 3'b000,
    SLL     = 3'b001,
    SLT     = 3'b010,
    SLTU    = 3'b011,
    XOR     = 3'b100,
    SRL_SRA = 3'b101,
    OR      = 3'b110,
    AND     = 3'b111
  } r_funct3_e;

  typedef enum logic [2:0] {
    ADDI      = 3'b000,
    SLLI      = 3'b001,
    SLTI      = 3'b010,
    SLTIU     = 3'b011,
    XORI      = 3'b100,
    SRLI_SRAI = 3'b101,
    ORI       = 3'b110,
    ANDI      = 3'b111
  } i_funct3_e;


  typedef enum logic [2:0] {
    SB = 3'b000,
    SH = 3'b001,
    SW = 3'b010
  } s_funct3_e;

  typedef enum logic [2:0] {
    LB  = 3'b000,
    LH  = 3'b001,
    LW  = 3'b010,
    LBU = 3'b100,
    LHU = 3'b101
  } l_funct3_e;

  typedef enum logic [2:0] {
    BEQ  = 3'b000,
    BNE  = 3'b001,
    BLT  = 3'b100,
    BGE  = 3'b101,
    BLTU = 3'b110,
    BGEU = 3'b111
  } b_funct3_e;

  typedef enum logic [2:0] {JALR = 3'b000} j_funct3_e;

  typedef enum logic [7:0] {
    SUB_SRA = 7'b0100000,
    OTHER   = 7'b0000000
  } r_funct7_e;

  typedef enum logic [7:0] {
    SRAI  = 7'b0100000,
    OTHER = 7'b0000000
  } i_funct7_e;

endpackage
