package package_uvm;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "mul_sequence_item.svh"
    `include "mul_sequence.svh"
    `include "mul_coverage_collector.svh"
    `include "mul_monitor.svh"
    `include "mul_driver.svh"
    `include "mul_agent.svh"
    `include "mul_scoreboard.svh"
    `include "mul_env.svh"
    `include "mul_test.svh"
endpackage : package_uvm