package package_uvm;
    import uvm_pkg::*;
     `include "uvm_macros.svh"
     //`include "riscv_pkg.sv"
     `include "alu_sequence_item.svh"
     `include "alu_sequence.svh"
     `include "alu_monitor.svh"
     `include "alu_driver.svh"
     `include "alu_sequencer.svh"
     `include "alu_agent.svh"
     `include "alu_scoreboard.svh"
     `include "alu_env.svh"
     `include "alu_test.svh"
endpackage : package_uvm