package package_uvm;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "riscv_pkg.sv"
    `include "scoreboard.svh"
    `include "subscriber.svh"
    `include "env.svh"
    `include "test.svh"
endpackage : package_uvm