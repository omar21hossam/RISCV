/*package riscv_classes_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "riscv_fetch_config_obj.svh"
    `include "riscv_seqitem.svh"
    `include "riscv_sequence_b.svh"
    `include "riscv_sequencer.svh"
    `include "riscv_main_driver.svh"
    `include "fetch_monitor.svh"
    `include "fetch_agent.svh"
    `include "riscv_scoreboard.svh"
    `include "riscv_subscriber.svh"
    `include "riscv_env.svh"
    `include "riscv_test.svh"
endpackage : riscv_classes_pkg*/
package riscv_classes_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"  
  `include "prefetch/riscv_config_obj.svh"
  `include "prefetch/riscv_seqitem.svh"
  `include "prefetch/fetch_seq_item.svh"
  `include "prefetch/riscv_sequence_b.svh"
  `include "prefetch/riscv_sequencer.svh"
  `include "prefetch/riscv_main_driver.svh"
  `include "prefetch/fetch_monitor.svh"
  `include "prefetch/fetch_agent.svh"
  `include "prefetch/fetch_scoreboard.svh"
  `include "prefetch/riscv_subscriber.svh"
  `include "riscv_env.svh"
  `include "riscv_test.svh"
endpackage