class lsu_sequence extends uvm_sequence;
  //==================================================================================
  // Registeration
  //==================================================================================
  `uvm_object_utils(lsu_sequence)

  //==================================================================================
  // Classes Handles
  //==================================================================================
  lsu_sequence_item m_seq_item;

  //==================================================================================
  // Function: Constructor
  //==================================================================================
  function new(string name = "lsu_sequence");
    super.new(name);
  endfunction

  //==================================================================================
  // Task: Pre-body
  //==================================================================================
  task pre_body();
    m_seq_item = lsu_sequence_item::type_id::create("m_seq_item");
  endtask

  //==================================================================================
  // Task: Body
  //==================================================================================
  task body();
    repeat (10000) begin
      start_item(m_seq_item);
      if (!m_seq_item.randomize())
        `uvm_fatal(get_name(), "Failed to randomize sequence item");
      finish_item(m_seq_item);
    end
  endtask

endclass
