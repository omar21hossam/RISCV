interface interface_clk (
    input logic clk
);

    logic monitor_done;  
endinterface